**inv**
* SPICE3 file created from inv.ext - technology: sky130A

.option scale=0.01u

.include ./pshort.lib
.include ./nshort.lib

//.subckt inv A Y VPWR VGND
M0 Y A VGND VGND nshort_model.0 ad=1435 pd=152 as=1365 ps=148 w=35 l=23  
M1 Y A VPWR VPWR pshort_model.0 ad=1443 pd=152 as=1517 ps=156 w=37 l=23

C0 A y 0.06fF
C1 Y VPWR 0.12fF
C2 A VPWR 0.27fF
C3 Y VGND 0.15fF
C4 A VGND 0.24fF
C5 VPWR VGND 0.49fF

* power sources excitation etc.
* v_instance_name posive_node negetive_node value
VDD VPWR 0 3.3V
VSS VGND 0 0
Va A GND PULSE(0 3.3 0 0.1n 0.1n 2n 4n)

.control
tran 1n 20n
setplot tran1
plot -VDD#branch
plot A Y
.endc
.end
