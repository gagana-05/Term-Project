* SPICE3 file created from inv.ext - technology: sky130A

.option scale=0.01u

.include ./pshort.lib
.include ./nshort.lib

.subckt inv A Y VPWR VGND
X0 Y A VGND VGND nshort_model.0 ad=1435 pd=152 as=1365 ps=148 w=35 l=23
X1 Y A VPWR VPWR pshort_model.0 ad=1443 pd=152 as=1517 ps=156 w=37 l=23
C0 A Y 0.06fF
C1 Y VPWR 0.12fF
C2 A VPWR 0.27fF
C3 Y VGND 0.15fF
C4 A VGND 0.24fF
C5 VPWR VGND 0.49fF
.ends

* power sources excitation etc.
* v_instance_name posive_node negetive_node value
VDD VPWR 0 3.3V
VSS VGND 0 0
Va A VGND PULSE(0V 3.3V 0 0.1ns 0.1ns 2ns 4ns)
.tran 1n 20n
.control
run
.endc
.end
